`timescale 1ns / 1ps

module TB_Shidt_Rows(  );

reg [127:0] shift_rows_in;
wire  [127:0] shift_row_out;

Shift_Rows S_R (shift_rows_in,shift_row_out);

initial 
begin
	$monitor("input= %H , output= %h",shift_rows_in,shift_row_out);
	shift_rows_in = 128'h_01020304_05060708_09101112_13141516;
	#10;
	shift_rows_in = 128'h_49ded289_45db96f1_7f39871a_7702533b;
	#10;
	shift_rows_in = 128'h_ac73cf7b_efc111df_13b5d6b5_45235ab8;
end

endmodule
