`timescale 1ns / 1ps

module TB_invarse_Shift_Rows(  );

reg [127:0] inv_shift_rows_in;
wire  [127:0] inv_shift_row_out;

inverse_shift_rows I_S_R1 (inv_shift_rows_in,inv_shift_row_out);

initial 
begin
	$monitor("input= %H , output= %h",inv_shift_rows_in,inv_shift_row_out);
	inv_shift_rows_in = 128'h01020304_05060708_09101112_13141516;
	#10;
	inv_shift_rows_in = 128'h338b762051667d92798febc20a3fbe67;
	#10;
	inv_shift_rows_in = 128'hac73cf7b_efc111df_13b5d6b5_45235ab8;
end

endmodule